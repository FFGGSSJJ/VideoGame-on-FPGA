//-------------------------------------------------------------------------
//    Ball.sv                                                            --
//    Viral Mehta                                                        --
//    Spring 2005                                                        --
//                                                                       --
//    Modified by Stephen Kempf 03-01-2006                               --
//                              03-12-2007                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Modified by Po-Han Huang  12-08-2017                               --
//    Spring 2018 Distribution                                           --
//                                                                       --
//    For use with ECE 385 Lab 8                                         --
//    UIUC ECE Department                                                --
//-------------------------------------------------------------------------


module  ball ( input         Clk,                // 50 MHz clock
                             Reset,              // Active-high reset signal
                             frame_clk,          // The clock indicating a new frame (~60Hz)
               input [9:0]   DrawX, DrawY,       // Current pixel coordinates
					input [7:0]	  keycode,
					input 		  collision,
               output logic  is_ball,             // Whether current pixel belongs to ball or background
					output logic [9:0]  Ball_X_Pos_out, Ball_Y_Pos_out, Ball_Size_out, Ball_Y_Step_out
              );
    
    parameter [9:0] Ball_X_Center = 10'd320;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center = 10'd240;  // Center position on the Y axis
    parameter [9:0] Ball_X_Min = 10'd0;       // Leftmost point on the X axis
    parameter [9:0] Ball_X_Max = 10'd639;     // Rightmost point on the X axis
    parameter [9:0] Ball_Y_Min = 10'd0;       // Topmost point on the Y axis
    parameter [9:0] Ball_Y_Max = 10'd479;     // Bottommost point on the Y axis
    parameter [9:0] Ball_Size = 10'd10;        // Ball size
    
    logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion;
    logic [9:0] Ball_X_Pos_in, Ball_X_Motion_in, Ball_Y_Pos_in, Ball_Y_Motion_in;
    logic [9:0] Ball_X_Step;      // Step size on the X axis
    logic [9:0] Ball_Y_Step;      // Step size on the Y axis	 
	 logic [9:0] counter;
	 
	 //output 
	 assign Ball_X_Pos_out = Ball_X_Pos;
	 assign Ball_Y_Pos_out = Ball_Y_Pos;
	 assign Ball_Size_out = Ball_Size;
	 assign Ball_Y_Step_out = Ball_Y_Step;
	 
	 
    //////// Do not modify the always_ff blocks. ////////
    // Detect rising edge of frame_clk
    logic frame_clk_delayed, frame_clk_rising_edge;
    always_ff @ (posedge Clk) begin
        frame_clk_delayed <= frame_clk;
        frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
    end
    // Update registers
    always_ff @ (posedge Clk)
    begin
        if (Reset)
        begin
            Ball_X_Pos <= Ball_X_Center;
            Ball_Y_Pos <= Ball_Y_Center;
				Ball_X_Step <= 10'd0;
				Ball_Y_Step <= 10'd0;
            Ball_X_Motion <= Ball_X_Step;
            Ball_Y_Motion <= Ball_Y_Step;
        end
        else
        begin
            Ball_X_Pos <= Ball_X_Pos_in;
            Ball_Y_Pos <= Ball_Y_Pos_in;
            Ball_X_Motion <= Ball_X_Motion_in;
            Ball_Y_Motion <= Ball_Y_Motion_in;
				if (frame_clk_rising_edge)
				begin
					if( Ball_Y_Pos + Ball_Size >= Ball_Y_Max )  // Ball is at the bottom edge, BOUNCE!
						 Ball_Y_Step <= ~10'd7+1;
					else if( Ball_X_Pos >= Ball_X_Max)  // Ball is at the right edge, BOUNCE!
						begin 
							Ball_X_Pos <= Ball_X_Pos_in + ~Ball_X_Max + 1'b1;
						end
					else if ( Ball_X_Pos <= Ball_X_Min)  // Ball is at the left edge, BOUNCE!
						begin
							Ball_X_Pos <= Ball_X_Pos_in + Ball_X_Max;
						end
					else if (collision == 1'b1)
						begin
							Ball_Y_Step <= ~10'd7+1;
						end
					else
						begin
							case(keycode)
								//Left
								8'h04: begin
											Ball_X_Step <= ~10'd1+1;
										end
								//Right
								8'h07: begin
											Ball_X_Step <= 10'd1;
										end
								default:
										begin
											Ball_X_Step <= 10'b0;
										end
							endcase
						end
						
						counter <= counter + 1'b1;
						if (counter>3)
						begin
							Ball_Y_Step <= Ball_Y_Step + 1'b1;
							counter <= 1'b0;
						end

				end
				
        end
    end
    //////// Do not modify the always_ff blocks. ////////
    
    // You need to modify always_comb block.
    always_comb
    begin
        // By default, keep motion and position unchanged
        Ball_X_Pos_in = Ball_X_Pos;
        Ball_Y_Pos_in = Ball_Y_Pos;
        Ball_X_Motion_in = Ball_X_Motion;
        Ball_Y_Motion_in = Ball_Y_Motion;
        
        // Update position and motion only at rising edge of frame clock
        if (frame_clk_rising_edge)
        begin
				Ball_X_Motion_in = Ball_X_Step;
				Ball_Y_Motion_in = Ball_Y_Step;
            Ball_X_Pos_in = Ball_X_Pos + Ball_X_Motion;
            Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;
        end
   
    end
    
    // Compute whether the pixel corresponds to ball or background
    /* Since the multiplicants are required to be signed, we have to first cast them
       from logic to int (signed by default) before they are multiplied. */
    int DistX1, DistY1, DistX2, DistY2, Size;
    assign DistX1 = DrawX - Ball_X_Pos;
    assign DistY1 = DrawY - Ball_Y_Pos;
    assign DistX2 = DrawX - Ball_X_Pos + Ball_X_Max;
    assign DistY2 = DrawY - Ball_Y_Pos;
    assign Size = Ball_Size;
    always_comb 
	 begin
        if (((DistX1*DistX1 + DistY1*DistY1) <= (Size*Size)) || ((DistX2*DistX2 + DistY2*DistY2) <= (Size*Size)))
            is_ball = 1'b1;
        else
            is_ball = 1'b0;
        /* The ball's (pixelated) circle is generated using the standard circle formula.  Note that while 
           the single line is quite powerful descriptively, it causes the synthesis tool to use up three
           of the 12 available multipliers on the chip! */
    end
    
endmodule
